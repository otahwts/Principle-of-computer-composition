LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY decoder0000 IS
    PORT (
        OP  : IN  STD_LOGIC_VECTOR(2 DOWNTO 0);
		  S  : OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
		 
);
END decoder0000;

ARCHITECTURE behav OF decoder0000 IS


BEGIN
		PROCESS(OP)
			BEGIN
				S <= '0'&OP;
			END PROCESS;

END behav;